


module params();

parameter data_bus_size = 16;
parameter addr_bus_size = 16;

endmodule
